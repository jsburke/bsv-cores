../../../Flute/src_Core/CPU/EX_ALU_functions.bsv