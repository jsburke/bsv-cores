../../../upstream/Flute/src_Core/CPU/IntMulDiv.bsv