../../../upstream/Flute/src_Core/CPU/CPU_Fetch_C.bsv