../../../Flute/src_Core/CPU/CPU_StageF.bsv