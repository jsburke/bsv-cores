../../../upstream/Flute/src_Core/CPU/CPU_StageD.bsv