../../../Flute/src_Core/CPU/RISCV_MBox.bsv