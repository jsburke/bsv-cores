../../../upstream/Flute/src_Core/CPU/CPU_Stage3.bsv