../../../upstream/Flute/src_Core/CPU/FBox_Top.bsv