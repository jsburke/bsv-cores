../../../upstream/Flute/src_Core/CPU/FBox_Core.bsv