../../../Flute/src_Core/CPU/CPU_IFC.bsv