../../../upstream/Flute/src_Core/CPU/CPU_Globals.bsv