../../../Flute/src_Core/CPU/Branch_Predictor.bsv