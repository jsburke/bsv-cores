../../../Flute/src_Core/CPU/CPU_Stage2.bsv