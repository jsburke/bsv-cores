../../../upstream/Flute/src_Core/CPU/FPU.bsv