../../../Flute/src_Core/CPU/CPU.bsv