../../../upstream/Flute/src_Core/CPU/Shifter_Box.bsv