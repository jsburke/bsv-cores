../../../Flute/src_Core/CPU/CPU_Decode_C.bsv