../../../upstream/Piccolo/src_Core/CPU/CPU.bsv