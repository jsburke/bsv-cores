../../../upstream/Flute/src_Core/CPU/CPU_Stage1.bsv